ONE-TRANSISTOR CIRCUIT (Fig. 1.2)
*
Q1 2 1 0 QMOD
RC 2 3 1K
RB 3 1 200K
VCC 3 0 5
*
.MODEL QMOD NPN IS=1E-16 BF=100
*
.OP
.END
